
module mystery_module (
    input a,
    input b,
    input c,
    output y
);

    assign y = a | c;

endmodule
