`timescale 1ns/1ps

module example2 (
    
);

    // reg / wire declarations here


endmodule
